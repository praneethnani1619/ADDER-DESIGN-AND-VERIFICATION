interface add_if;
  logic clk;
  logic reset;
  logic [7:0] ip1;   
  logic [7:0] ip2;   
  logic [8:0] out;
endinterface
